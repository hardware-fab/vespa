//----------------------------------------------------------------------------
//  This file is a part of the VESPA SoC Prototyping Framework
//
//  This program is free software; you can redistribute it and/or modify
//  it under the terms of the Apache 2.0 License.
//
// File:    bram18.py
// Authors: Gabriele Montanaro
//          Andrea Galimberti
//          Davide Zoni
// Company: Politecnico di Milano
// Mail:    name.surname@polimi.it
//
//----------------------------------------------------------------------------

module bram18 #(  
    parameter READ_WIDTH            = 18,
    parameter WRITE_WIDTH           = 18,
    parameter ADDR_WIDTH            = 10,
    parameter WE_WIDTH              = 2
    )
    (
    input                        clk,
    input                        reset,
    input  [ADDR_WIDTH-1:0]      addr_i,
    input                        valid_i,
    output [READ_WIDTH-1:0]      data_o
    );
    wire [WRITE_WIDTH-1:0] data_i ;
    wire [WE_WIDTH-1:0]    we ;
    wire                   regce;
    assign  we      = { WE_WIDTH{1'b0}    };
    assign  data_i  = { WRITE_WIDTH{1'b0} };
    assign  regce   = 1'b0;
    BRAM_SINGLE_MACRO #(
        .BRAM_SIZE("18Kb"), // Target BRAM, "18Kb" or "36Kb" 
        .DEVICE("7SERIES"), // Target Device: "7SERIES" 
        .DO_REG(0), // Optional output register (0 or 1)
        .INIT(18'b000000000000000000), // Initial values on output port
        .INIT_FILE ("NONE"),
        .WRITE_WIDTH(WRITE_WIDTH), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .READ_WIDTH(READ_WIDTH),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .SRVAL(18'b000000000000000000), // Set/Reset value for port output
        .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        .INIT_00(256'h28002500230020001e001b0019001600140011000f000c000a00070005000200),
.INIT_01(256'h32003200320032003200320032003200320032003200320032002f002d002a00),
.INIT_02(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_03(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_04(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_05(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_06(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_07(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_08(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_09(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_0A(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_0B(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_0C(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_0D(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_0E(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_0F(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_10(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_11(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_12(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_13(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_14(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_15(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_16(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_17(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_18(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_19(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1A(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1B(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1C(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1D(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1E(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1F(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_20(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_21(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_22(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_23(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_24(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_25(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_26(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_27(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_28(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_29(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2A(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2B(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2C(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2D(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2E(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2F(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_30(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_31(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_32(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_33(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_34(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_35(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_36(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_37(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_38(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_39(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3A(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3B(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3C(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3D(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3E(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3F(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INITP_00(256'h0000000000000000000000000000000000000000000000000000001111111111),
.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)) 
        BRAM_SINGLE_MACRO_inst (
            .DO(data_o),   // Output data, width defined by READ_WIDTH parameter
            .ADDR(addr_i), // Input address, width defined by read/write port depth look at the table below
            .CLK(clk),     // 1-bit input clock
            .DI(data_i),   // Input data port, width defined by WRITE_WIDTH parameter
            .EN(valid_i),  // 1-bit input RAM enable
            .REGCE(regce), // 1-bit input output register enable
            .RST(reset),   // 1-bit input reset
            .WE(we)        // Input write enable, width defined by write port depth look at tabel below
        );
        /////////////////////////////////////////////////////////////////////
        //  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            //
        // WRITE_WIDTH |           | WRITE Depth |            |  WE Width  //
        // ============|===========|=============|============|============//
        //    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   //
        //    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   //
        //    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   //
        //    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   //
        //    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   //
        //     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   //
        //     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   //
        //     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   //
        //     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   //
        //       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   //
        //       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   //
        //       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   //
        //       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   //
        /////////////////////////////////////////////////////////////////////
        
 endmodule